//assign 连续赋值语句是把右边赋值给左边，assign left_side = right_side;
module top_module(
    input in,
    output out
);

assign out = in;

endmodule