module top_modle (
    output zero
);

endmodule


module top_modle (
    zero
);
  output zero;
endmodule
//两种方式都可以构建一个没有输入，只有输出，并且输出为0的电路