module top_module (
    input  a,
    b,
    c,
    output w,
    x,
    y,
    z
);

  assign w = a;
  assign x = b;
  assign y = c;
  assign z = d;


endmodule
//{'a,b,c,d'}注意逗号的使用